module data_mem
(
    input clock
);

endmodule