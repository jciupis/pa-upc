module data_mem
(
    input clock,
    input read_cmd,
    input write_cmd,
    input byte_access,
    input  [31:0] address,
    output [31:0] data
);

endmodule